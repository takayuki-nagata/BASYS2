library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity SSegDecoder is
	Port (
		DIG :  in std_logic_vector (3 downto 0);
		LED : out std_logic_vector (6 downto 0)
	);
end SSegDecoder;

architecture Behavioral of SSegDecoder is
begin
	process(DIG) begin
		case DIG is
			when "0000" => LED <= "0000001"; -- 0
			when "0001" => LED <= "1001111"; -- 1
			when "0010" => LED <= "0010010"; -- 2
			when "0011" => LED <= "0000110"; -- 3
			when "0100" => LED <= "1001100"; -- 4
			when "0101" => LED <= "0100100"; -- 5
			when "0110" => LED <= "0100000"; -- 6
			when "0111" => LED <= "0001111"; -- 7
			when "1000" => LED <= "0000000"; -- 8
			when "1001" => LED <= "0000100"; -- 9
			when others => LED <= "XXXXXXX";
		end case;
	end process;
end Behavioral;